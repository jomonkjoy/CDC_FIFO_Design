module cpu_if_cdc (
);

endmodule
